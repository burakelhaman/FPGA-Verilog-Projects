module grayverilog(input x,clk,h, output reg[6:0]disp);
reg[3:0]count=0;
always@(posedge clk)begin
	if (h==0)begin
		if (x==1) count=count+1;
		
		else		count=count-1;
	end
	
case (count)
	4'b0000:disp = 7'b1111110;
	4'b0001:disp = 7'b0110000;
	4'b0010:disp = 7'b1101101;
	4'b0011:disp = 7'b1111001;
	4'b0100:disp = 7'b0110011;
	4'b0101:disp = 7'b1011011;
	4'b0110:disp = 7'b1011111;
	4'b0111:disp = 7'b1110000;
	4'b1000:disp = 7'b1111111;
	4'b1001:disp = 7'b1111011;
	4'b1010:disp = 7'b1111101;
	4'b1011:disp = 7'b0011111;
	4'b1100:disp = 7'b1001110;
	4'b1101:disp = 7'b0111101;
	4'b1110:disp = 7'b1001111;
	4'b1111:disp = 7'b1000111;
endcase
end
endmodule
